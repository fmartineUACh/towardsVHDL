library verilog;
use verilog.vl_types.all;
entity cy_6gserdes_core is
    port(
        txda            : in     vl_logic_vector(7 downto 0);
        txdb            : in     vl_logic_vector(7 downto 0);
        txdc            : in     vl_logic_vector(7 downto 0);
        txdd            : in     vl_logic_vector(7 downto 0);
        txpera          : out    vl_logic;
        txperb          : out    vl_logic;
        txperc          : out    vl_logic;
        txperd          : out    vl_logic;
        txcta           : in     vl_logic_vector(1 downto 0);
        txctb           : in     vl_logic_vector(1 downto 0);
        txctc           : in     vl_logic_vector(1 downto 0);
        txctd           : in     vl_logic_vector(1 downto 0);
        txopa           : in     vl_logic;
        txopb           : in     vl_logic;
        txopc           : in     vl_logic;
        txopd           : in     vl_logic;
        txclka          : in     vl_logic;
        txclkb          : in     vl_logic;
        txclkc          : in     vl_logic;
        txclkd          : in     vl_logic;
        txclko          : out    vl_logic;
        txrate          : in     vl_logic;
        txmode          : in     vl_logic_vector(1 downto 0);
        txcksel         : in     vl_logic;
        txrstb          : in     vl_logic;
        scsel           : in     vl_logic;
        rxda            : out    vl_logic_vector(7 downto 0);
        rxdb            : out    vl_logic_vector(7 downto 0);
        rxdc            : out    vl_logic_vector(7 downto 0);
        rxdd            : out    vl_logic_vector(7 downto 0);
        rxsta           : out    vl_logic_vector(2 downto 0);
        rxstb           : out    vl_logic_vector(2 downto 0);
        rxstc           : out    vl_logic_vector(2 downto 0);
        rxstd           : out    vl_logic_vector(2 downto 0);
        rxopa           : out    vl_logic;
        rxopb           : out    vl_logic;
        rxopc           : out    vl_logic;
        rxopd           : out    vl_logic;
        rxrate          : in     vl_logic;
        rfen            : in     vl_logic;
        rxmode          : in     vl_logic_vector(1 downto 0);
        rxcksel         : in     vl_logic;
        framchar        : in     vl_logic;
        rfmode          : in     vl_logic;
        decmode         : in     vl_logic;
        parctl          : in     vl_logic;
        spdsel          : in     vl_logic;
        rxclka          : out    vl_logic;
        rxclkb          : inout  vl_logic;
        rxclkc          : out    vl_logic;
        rxclkd          : inout  vl_logic;
        lesstime        : in     vl_logic;
        resetb          : out    vl_logic;
        refclk          : in     vl_logic;
        warning_disable : in     vl_logic;
        serial_outa1    : out    vl_logic;
        serial_outb1    : out    vl_logic;
        serial_outc1    : out    vl_logic;
        serial_outd1    : out    vl_logic;
        serial_outa2    : out    vl_logic;
        serial_outb2    : out    vl_logic;
        serial_outc2    : out    vl_logic;
        serial_outd2    : out    vl_logic;
        serial_ina1     : in     vl_logic;
        serial_inb1     : in     vl_logic;
        serial_inc1     : in     vl_logic;
        serial_ind1     : in     vl_logic;
        serial_ina2     : in     vl_logic;
        serial_inb2     : in     vl_logic;
        serial_inc2     : in     vl_logic;
        serial_ind2     : in     vl_logic;
        insela          : in     vl_logic;
        inselb          : in     vl_logic;
        inselc          : in     vl_logic;
        inseld          : in     vl_logic;
        sdasel          : in     vl_logic;
        lpen            : in     vl_logic;
        oele            : in     vl_logic;
        bistle          : in     vl_logic;
        rxle            : in     vl_logic;
        boe             : in     vl_logic_vector(7 downto 0);
        bondst          : inout  vl_logic_vector(1 downto 0);
        masterb         : in     vl_logic;
        bond_all        : inout  vl_logic;
        bond_inhb       : in     vl_logic;
        lfiab           : out    vl_logic;
        lfibb           : out    vl_logic;
        lficb           : out    vl_logic;
        lfidb           : out    vl_logic;
        trstzb          : in     vl_logic;
        recovered_clka  : out    vl_logic;
        recovered_clkb  : out    vl_logic;
        recovered_clkc  : out    vl_logic;
        recovered_clkd  : out    vl_logic;
        clkadj_a        : out    vl_logic;
        clkadj_b        : out    vl_logic;
        clkadj_c        : out    vl_logic;
        clkadj_d        : out    vl_logic;
        out1pwrdn       : out    vl_logic_vector(3 downto 0);
        out2pwrdn       : out    vl_logic_vector(3 downto 0)
    );
end cy_6gserdes_core;
