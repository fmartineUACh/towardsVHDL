
package VERIBEST is

    --  Reserved for future use

end package VERIBEST;


