--	This design describes a simple SERDES application for a PSI device that transmits 
--	the 16-bit output of four side-by-side 4-bit counters and resets or channels the received
-- data to be presented at the PSI outputs.
--	The 4-bit counters are incremented at every transmit clock cycle and wraps around to 
--	"0000" after reaching the maximum count value of "1111".  When a line fault is 
--	detected on the receiver, the SERDES output signal lfib is set to '0' and the data 
--	sequence "1111111100000000" is transmitted instead of the counter outputs.  
-- On the receive side, the design input signal "reset_rxd" controls whether the received 
-- data bits are reset.  When reset_rxd is '1', all 16-bits of received data are set to '0'.  
--	Otherwise, it is left as is.  Also, when test mode is enabled (test_en = '1'), both 
--	line loopback and diagnostic loopback are enabled.  The user may also specify these 
--	two loopback modes externally through the "lineloop_en" and "diagloop_en" input ports. 


library ieee;
use ieee.std_logic_1164.all;
library cypress;
use cypress.rtlpkg.all;
use cypress.std_arith.all;

entity PSI is port(  
	 -- reference differential clock
	 refclk_p, refclk_n: in std_logic;   	
	 -- serial differential input
	 serial_inn, serial_inp: in std_logic;  
	 -- signal detect
	 sd: in std_logic;
	 -- synchronous reset for 16-bit receive data 						
	 reset_rxd:  in std_logic;
	 -- control signal, enables test mode					
	 test_en: in std_logic;
	 -- enables line loop on serial transmit data 			    
	 lineloop_en:  in std_logic;
	 -- enables diagnostic loopback of transmit data	
	 diagloop_en:  in std_logic;
	 -- Lock to Reference clock select
	 lockrefb: in std_logic;
	 -- FIFO reset
	 fifo_rstb: in std_logic;
	 -- Loop Timing mode select
	 loop_time: in std_logic;
	 -- line loopback mode (non-retimed data) enable
	 loopa: in std_logic;
	 -- all logic circuit reset
  	 resetb: in std_logic;
	 -- Power down enable
	 pwrdnb: in std_logic;
	 -- FIFO error status
	 fifo_err: out std_logic;
	 -- serial differential output
	 serial_outn, serial_outp: out std_logic;
	 -- 16-bit receive data output to pins
	 rxdata_out: out std_logic_vector (15 downto 0) 
	
);
end PSI;

architecture PSI_arch of PSI is

	-- 16-bit transmit data generated by counters in macrocell register
	signal txdata: std_logic_vector (15 downto 0);
	-- 16-bit transmit data registered output to SERDES	
 	signal txdata_out: std_logic_vector (15 downto 0);
	-- 16-bit receive data registered input from the SERDES
   signal rxdata_in: std_logic_vector (15 downto 0);
	-- 16-bit receive data input to macrocell register
	signal rxdata: std_logic_vector (15 downto 0);
	-- 16-bit processed receive data	output from macrocell register
	signal rxdata_reg: std_logic_vector (15 downto 0); 
	-- transmit and receive clocks
	signal txclk, rxclk: std_logic;
	-- diagloop control signal			
	signal diagloop_sel: std_logic;
	-- lineloop control signal			
	signal lineloop_sel: std_logic;
	-- line fault indicator signal			
	signal linedown:std_logic;		
	
	

begin

	-- instantiate the SERDES
	U1: cy_25g01serdes	
		port map(
			txd          => txdata_out,
			fifo_rstb    => fifo_rstb,			
			loop_time    => loop_time,		
			diagloop     => diagloop_sel,
			loopa        => loopa,			
			lineloop     => lineloop_sel,
			resetb       => resetb,		
			pwrdnb       => pwrdnb,			
			lockrefb     => lockrefb,		
			refclk_n     => refclk_n,
			refclk_p     => refclk_p,
			serial_in_n  => serial_inn,
			serial_in_p  => serial_inp,
			sd           => sd,
			serial_out_n => serial_outn,
			serial_out_p => serial_outp,
			fifo_err     => fifo_err,
			txclk        => txclk,
			rxd          => rxdata_in,
			rxclk        => rxclk,
			lfib         => linedown
		);

	-- process the diagloop and lineloop control signals
	lineloop_sel <= lineloop_en or test_en;
	diagloop_sel <= diagloop_en or test_en;
	
	-- Generate transmit data from counter output when rising transmit clock edge occurs
	process (txclk)
	begin
		if (txclk'event and txclk='1') then
			if (linedown = '0') then
				txdata <= "1111111100000000";
			else
				txdata(15 downto 12) <= txdata(15 downto 12) + 1;
			 	txdata(11 downto 8) <= txdata(11 downto 8) + 1;
				txdata(7 downto 4) <= txdata(7 downto 4) + 1;
			 	txdata(3 downto 0) <= txdata(3 downto 0) + 1;
			end if;
		end if;
	end process;

	-- register transmit data before output to SERDES
	process (txclk)
	begin
		if (txclk'event and txclk='1') then
			txdata_out <= txdata;
		end if;
	end process;

	-- register receive data input from SERDES
	process (rxclk)
	begin
		if (rxclk'event and rxclk='1') then
			rxdata <= rxdata_in;
		end if;
	end process;

	-- register and process receive data at a macrocell
	process (rxclk)
	begin
		if (rxclk'event and rxclk='1') then
			if (reset_rxd = '1') then
				rxdata_reg <= (others => '0');
			else
				rxdata_reg <= rxdata;
			end if;
		end if;
	end process;

	-- register processed receive data before output to PSI pins
	process (rxclk)
	begin
		if (rxclk'event and rxclk='1') then
			rxdata_out <= rxdata_reg;
		end if;
	end process;
end PSI_arch;
