LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SELECT1 IS
    PORT (SNICKERS : IN X01Z
        ; MARS : IN X01Z
        ; MOUNDS : IN X01Z
        ; HERSHEYS : IN X01Z
        ; ENABLE : IN X01Z
        ; SNICKERS_OUT : OUT X01Z
        ; MARS_OUT : OUT X01Z
        ; MOUNDS_OUT : OUT X01Z
        ; HERSHEYS_OUT : OUT X01Z
        ; SEL_MADE : OUT X01Z
);

END SELECT1;

ARCHITECTURE A1 OF SELECT1 IS

    ATTRIBUTE ENUM_TYPE_ENCODING: STRING;

    SIGNAL FB_SNICKERS_OUT : X01Z;
    SIGNAL FB_MARS_OUT : X01Z;
    SIGNAL FB_MOUNDS_OUT : X01Z;
    SIGNAL FB_HERSHEYS_OUT : X01Z;

BEGIN 
    SNICKERS_OUT <= FB_SNICKERS_OUT ;
    MARS_OUT <= FB_MARS_OUT ;
    MOUNDS_OUT <= FB_MOUNDS_OUT ;
    HERSHEYS_OUT <= FB_HERSHEYS_OUT ;
    FB_SNICKERS_OUT <= ((SNICKERS AND ENABLE));
    FB_MARS_OUT <= ((MARS AND ENABLE));
    FB_MOUNDS_OUT <= ((MOUNDS AND ENABLE));
    FB_HERSHEYS_OUT <= ((HERSHEYS AND ENABLE));
    SEL_MADE <= ((((FB_SNICKERS_OUT OR FB_MARS_OUT) OR FB_MOUNDS_OUT) OR FB_HERSHEYS_OUT));


END A1;
