--------------------------------------------------------------------------------
--
--  Copyright Cypress Semiconductor Corporation, 1995,1996
--  as an unpublished work.
--

--------------------------------------------------------------------------------

PACKAGE int_arith is

    -- This is a dummy package for the clause "use cypress.int_arith.all;".

end int_arith;
