package gatespkg is
component and2 port(a,b:in bit; q:out bit); end component;
component or2 port(a,b:in bit; q:out bit); end component;
component inv port(a:in bit; qn:out bit); end component;
end package;


